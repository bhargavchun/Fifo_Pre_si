package fifo_pkg;
    `include "trans_fifo.sv"
    `include "driv_fifo.sv"
    `include "gen_fifo.sv"
    `include "mon_fifo.sv"
    `include "scb_fifo.sv"
    
    `include "environment.sv"
    
endpackage
